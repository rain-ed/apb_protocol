import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../../uvm_apb/tb/uvm_seq_item.sv"
`include "../../uvm_apb/tb/uvm_seq.sv"
`include "../../uvm_apb/tb/uvm_sqr.sv"
`include "../../uvm_apb/tb/uvm_drv.sv"
`include "../../uvm_apb/tb/uvm_mon.sv"
`include "../../uvm_apb/tb/uvm_agent.sv"
`include "../../uvm_apb/tb/uvm_scb.sv"
`include "../../uvm_apb/tb/uvm_env.sv"
`include "../../uvm_apb/tb/uvm_test.sv"
`include "../../uvm_apb/tb/uvm_interface.sv"
`include "../../uvm_apb/tb/uvm_dut.sv"
`include "../../uvm_apb/tb/uvm_tb_top.sv"
